/****************************************************************************/
/**
 * \file <FILE_NAME>
 * 
 * \date <YYYY-MM-DD>
 * 
 * \author <YOUR_NAME>
 * 
 * \brief ...
 * 
 * \details ...
 * 
 * \see
 */
/****************************************************************************/

`ifndef _TEMPLATE_H
`define _TEMPLATE_H

`define timescale 1ns

`endif // _TEMPLATE_H
