/****************************************************************************/
/**
 * \file      timescale
 *
 * \project   -
 *
 * \langv     Verilog-2005
 *
 * \brief     Define the timescale.
 *
 * \details   Every Verilog module should contain the definition of the
 *            timescale directive, either by defining it or by including an
 *            apropriate header file like this one.
 *
 * \bug       -
 *
 * \see       -
 *
 * \copyright GPLv2
 *
 * Revision history:
 *
 * \version   0.1
 * \date      2015-06-04
 * \author    Andreas Mueller
 */
/****************************************************************************/

`ifndef timescale
`define timescale 1 ns / 1 ps
`endif
