/****************************************************************************/
/**
 * \file      timescale
 *
 * \project   -
 *
 * \langv     Verilog-2005
 *
 * \brief     Define the timescale.
 *
 * \details   Every Verilog module should contain the definition of the
 *            timescale directive, either by defining it or by including an
 *            appropriate header file like this one.
 *
 * \bug       -
 *
 * \see       -
 *
 * \copyright GPLv2
 *
 * Revision history:
 *
 * \version   0.1
 * \date      2015-06-04
 * \author    Andreas Mueller
 */
/****************************************************************************/

`ifndef _H_TIMESCALE
`timescale 10 ns / 1 ns
`endif // _H_TIMESCALE
