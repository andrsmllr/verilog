/**
 * \file      qsgmii.vh
 *
 * \project   mii_lib
 *
 * \langv     Verilog-2005
 *
 * \brief     Macros for the quad serial gigabit media-independent interface (QSGMII).
 *
 * \details   This file contains macros for the quad serial gigabit
 *            media-independent interface (QSGMII).
 *            These macros are intended as a uniform way to easily add QSGMIIs
 *            to the port interface of a module or to quickly declare nets of
 *            the required types.
 *
 * \bug      -
 *
 * \see      -
 *
 * \copyright GPLv2
 *
 * Revision history:
 *
 * \version   0.1
 * \date      2015-11-25
 * \author    Andreas Mueller
 * \brief     Create file.
**/

`ifndef _QSGMII_H
`define _QSGMII_H

/**
 * Quad serial gigabit media-independent interface (QSGMII).
**/
`define QSGMII(_type, _prefix, _suffix)
// This macro is a stub. TODO

`endif // _QSGMII_H
