/**
 * \file      <FILE_NAME>
 *
 * \project   <PROJECT_NAME>
 *
 * \langv     Verilog-2005
 *
 * \brief     <BRIEF_DESCRIPTION>
 *
 * \details   <DETAILED_DESCRIPTION>
 *
 * \bug       <BUGS_OR_KNOWN_ISSUES>
 *
 * \see       <REFERENCES>
 *
 * \copyright <COPYRIGHT_OR_LICENSE>
 *
 * Revision history:
 *
 * \version   <VERSION>
 * \date      <YYYY-MM-DD>
 * \author    <AUTHOR_NAME>
 * \brief     <BRIEF_DESCRIPTION>
**/

`ifndef _TEMPLATE_H
`define _TEMPLATE_H

`endif // _TEMPLATE_H

