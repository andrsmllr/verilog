/**
 * \file <FILE_NAME>
 * 
 * \date <YYYY-MM-DD>
 * 
 * \author <YOUR_NAME>
 * 
 * \brief ...
 * 
 * \details ...
 * 
 * \see
 */

/****************************************************************************/

module TESTBENCH_NAME
#(
    parameter PARAM1 = 0,
    parameter PARAM2 = 8
)
(
);


endmodule

