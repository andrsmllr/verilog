// Usually the modules to be instantiated reside in a different file wich must
// be included first.
`include "module_definition.v"

module module_instantiation;

// Verilog-1995 module instantiation.


// Verilog-2001 module instantiation.


// Verilog-2005 module instantiation.


endmodule
