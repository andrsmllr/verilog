module system_functions;

endmodule
