module system_tasks;

endmodule
