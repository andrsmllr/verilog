/**
 * \file      dvbc_qam_mapper_tb
 *
 * \project   dvbc
 *
 * \langv     Verilog-2005
 *
 * \brief     Testbench for QAM mapper for DVB-C modulator.
 *
 * \details   -
 *
 * \bug       -
 *
 * \see       -
 *
 * \copyright GPLv2
 *
 * Revision history:
 *
 * \version   0.1
 * \date      2015-06-05
 * \author    Andreas Mueller
**/

module dvbc_qam_mapper_tb
#(
    parameter PARAM1 = 0,
    parameter PARAM2 = 8
)
(
);


endmodule

