/**
 * \file      dvbc_qam_mapper_tb
 *
 * \project   dvbc
 *
 * \langv     Verilog-2005
 *
 * \brief     Testbench for QAM mapper for DVB-C modulator.
 *
 * \details   -
 *
 * \bug       -
 *
 * \see       -
 *
 * \copyright GPLv2
 *
 * Revision history:
 *
 * \version   0.1
 * \date      2015-06-05
 * \author    Andreas Mueller
 * \brief     Create file.
**/

module dvbc_qam_mapper_tb
#(
)
(
);

endmodule
