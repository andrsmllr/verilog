
`define PAD(signal, before, after) {{before'b0}, signal, {after'b0}}
`define TRIM(signal, left, right)

module pad_and_trim;

endmodule
