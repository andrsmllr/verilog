/**
 * \file      dvbc_randomizer_tb
 *
 * \project   dvbc
 *
 * \langv     Verilog-2005
 *
 * \brief     Testbench for randomizer to perform energy dispersal.
 *
 * \details   -
 *
 * \bug       -
 *
 * \see       -
 *
 * \copyright GPLv2
 *
 * Revision history:
 *
 * \version   0.1
 * \date      2015-06-05
 * \author    Andreas Mueller
**/

module dvbc_randomizer_tb
#(
    parameter PARAM1 = 0,
    parameter PARAM2 = 8
)
(
);


endmodule

